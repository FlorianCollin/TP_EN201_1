library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity trans is
    port (
        forward, play_pause, restart : in std_logic;
        nb_binaire : in std_logic_vector(9 downto 0); -- sortie de cpt_1_599
        nb_binaire_volume : in std_logic_vector(3 downto 0); --sortie de cpt_1_9
        s_cent, s_diz, s_unit : out std_logic_vector(6 downto 0);
        s_unit_vol : out std_logic_vector(6 downto 0);
        sortie1, sortie2, sortie3, sortie4 : out std_logic_vector(6 downto 0)
    );
end trans;

architecture behav of trans is

begin

    process(forward, play_pause, restart, nb_binaire, nb_binaire_volume)
    begin

        if (play_pause = '0') and (restart = '1') and (forward = '0') then
            -- Etat init
            sortie1 <= "0110001"; -- '['
            sortie2 <= "1111110"; -- '-'
            sortie3 <= "1111110"; -- '-'
            sortie4 <= "0000111"; -- ']'

        elsif (play_pause = '0') and (restart = '1') and (forward = '0') then
            -- Etat play fwd
            sortie1 <= "1111110"; -- '-'
            sortie2 <= "1111110"; -- '-'
            sortie3 <= "1111110"; -- '-'
            sortie4 <= "0000111"; -- ']'

        elsif (play_pause = '0') and (restart = '1') and (forward = '0') then
            -- Etat play bwd
            sortie1 <= "0110001"; -- '['
            sortie2 <= "1111110"; -- '-'
            sortie3 <= "1111110"; -- '-'
            sortie4 <= "1111110"; -- '-'

        elsif (play_pause = '0') and (restart = '1') and (forward = '0') then
            -- Etat pause
            sortie1 <= "1111110"; -- '-'
            sortie2 <= "1111110"; -- '-'
            sortie3 <= "1111110"; -- '-'
            sortie4 <= "1111110"; -- '-'

        elsif (play_pause = '0') and (restart = '1') and (forward = '0') then
            -- Etat stop
            sortie1 <= "0110001"; -- '['
            sortie2 <= "1111110"; -- '-'
            sortie3 <= "1111110"; -- '-'
            sortie4 <= "0000111"; -- ']'

        end if;

        case nb_binaire_volume is

            when "0001" => --1
                s_unit_vol <= "1001111";
            
            when "0010" =>
                s_unit_vol <= "0010010";
            
            when "0011" =>
                s_unit_vol <= "0000110";

            when "0100" =>
                s_unit_vol <= "1001100";
            
            when "0101" =>
                s_unit_vol <= "0100100"; 
            
            when "0110" =>
                s_unit_vol <= "0100000";
            
            when "0111" =>
                s_unit_vol <= "0001111";
            
            when "1000" =>
                s_unit_vol <= "0000000";
            
            when "1001" => -- 9
                s_unit_vol <= "0000100";

            when others =>
                s_unit_vol <= "0000100";

        end case;
            
        -- hihi ;)
        case (nb_binaire) is
            
            --when "0000000000" =>
                --s_unit <= "0000001";
                --s_diz <= "0000001";
                --s_cent <= "0000001";
            
            when "0000000001" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000010" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000011" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000100" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000101" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000110" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000000111" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000001000" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000001001" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "0000001010" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000001011" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000001100" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000001101" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000001110" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000001111" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000010000" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000010001" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000010010" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000010011" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "0000010100" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000010101" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000010110" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000010111" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011000" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011001" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011010" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011011" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011100" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011101" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "0000011110" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000011111" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100000" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100001" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100010" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100011" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100100" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100101" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100110" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000100111" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "0000101000" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101001" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101010" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101011" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101100" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101101" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101110" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000101111" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000110000" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000110001" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "0000110010" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000110011" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000110100" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000110101" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000110110" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000110111" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000111000" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000111001" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000111010" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000111011" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "0000111100" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0000111101" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0000111110" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0000111111" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000000" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000001" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000010" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000011" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000100" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000101" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "0001000110" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001000111" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001000" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001001" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001010" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001011" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001100" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001101" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001110" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001001111" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "0001010000" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010001" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010010" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010011" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010100" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010101" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010110" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001010111" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001011000" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001011001" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "0001011010" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001011011" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001011100" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001011101" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001011110" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001011111" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001100000" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001100001" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001100010" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001100011" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "0001100100" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001100101" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001100110" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001100111" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101000" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101001" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101010" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101011" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101100" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101101" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "0001101110" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001101111" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110000" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110001" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110010" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110011" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110100" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110101" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110110" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001110111" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "0001111000" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111001" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111010" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111011" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111100" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111101" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111110" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0001111111" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0010000000" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0010000001" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "0010000010" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010000011" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010000100" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010000101" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010000110" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010000111" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010001000" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010001001" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010001010" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010001011" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "0010001100" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010001101" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010001110" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010001111" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010000" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010001" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010010" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010011" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010100" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010101" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "0010010110" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010010111" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011000" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011001" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011010" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011011" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011100" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011101" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011110" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010011111" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "0010100000" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100001" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100010" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100011" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100100" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100101" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100110" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010100111" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010101000" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010101001" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "0010101010" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010101011" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010101100" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010101101" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010101110" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010101111" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010110000" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010110001" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010110010" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010110011" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "0010110100" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010110101" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010110110" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010110111" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111000" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111001" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111010" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111011" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111100" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111101" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "0010111110" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0010111111" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000000" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000001" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000010" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000011" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000100" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000101" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000110" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011000111" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "0011001000" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001001" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001010" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001011" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001100" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001101" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001110" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011001111" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011010000" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011010001" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "0011010010" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011010011" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011010100" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011010101" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011010110" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011010111" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011011000" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011011001" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011011010" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011011011" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "0011011100" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011011101" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011011110" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011011111" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100000" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100001" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100010" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100011" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100100" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100101" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "0011100110" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011100111" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101000" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101001" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101010" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101011" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101100" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101101" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101110" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011101111" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "0011110000" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110001" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110010" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110011" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110100" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110101" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110110" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011110111" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011111000" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011111001" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "0011111010" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0011111011" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0011111100" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0011111101" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0011111110" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0011111111" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0100000000" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0100000001" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0100000010" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0100000011" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "0100000100" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100000101" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100000110" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100000111" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001000" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001001" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001010" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001011" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001100" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001101" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "0010010";
            
            when "0100001110" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100001111" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010000" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010001" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010010" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010011" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010100" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010101" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010110" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100010111" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "0010010";
            
            when "0100011000" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011001" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011010" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011011" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011100" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011101" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011110" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100011111" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100100000" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100100001" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "0010010";
            
            when "0100100010" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100100011" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100100100" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100100101" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100100110" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100100111" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100101000" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100101001" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100101010" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100101011" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0010010";
            
            when "0100101100" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100101101" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100101110" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100101111" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110000" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110001" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110010" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110011" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110100" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110101" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0000110";
            
            when "0100110110" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100110111" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111000" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111001" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111010" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111011" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111100" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111101" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111110" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0100111111" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0000110";
            
            when "0101000000" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000001" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000010" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000011" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000100" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000101" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000110" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101000111" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101001000" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101001001" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0000110";
            
            when "0101001010" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101001011" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101001100" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101001101" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101001110" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101001111" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101010000" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101010001" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101010010" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101010011" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0000110";
            
            when "0101010100" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101010101" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101010110" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101010111" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011000" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011001" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011010" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011011" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011100" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011101" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0000110";
            
            when "0101011110" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101011111" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100000" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100001" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100010" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100011" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100100" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100101" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100110" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101100111" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "0000110";
            
            when "0101101000" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101001" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101010" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101011" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101100" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101101" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101110" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101101111" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101110000" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101110001" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "0000110";
            
            when "0101110010" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101110011" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101110100" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101110101" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101110110" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101110111" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101111000" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101111001" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101111010" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101111011" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "0000110";
            
            when "0101111100" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0101111101" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0101111110" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0101111111" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000000" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000001" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000010" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000011" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000100" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000101" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "0000110";
            
            when "0110000110" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110000111" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001000" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001001" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001010" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001011" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001100" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001101" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001110" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110001111" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0000110";
            
            when "0110010000" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010001" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010010" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010011" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010100" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010101" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010110" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110010111" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110011000" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110011001" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "1001100";
            
            when "0110011010" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110011011" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110011100" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110011101" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110011110" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110011111" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110100000" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110100001" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110100010" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110100011" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "1001100";
            
            when "0110100100" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110100101" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110100110" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110100111" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101000" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101001" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101010" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101011" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101100" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101101" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "1001100";
            
            when "0110101110" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110101111" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110000" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110001" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110010" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110011" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110100" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110101" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110110" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110110111" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "1001100";
            
            when "0110111000" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111001" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111010" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111011" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111100" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111101" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111110" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0110111111" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0111000000" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0111000001" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "1001100";
            
            when "0111000010" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111000011" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111000100" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111000101" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111000110" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111000111" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111001000" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111001001" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111001010" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111001011" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "1001100";
            
            when "0111001100" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111001101" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111001110" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111001111" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010000" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010001" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010010" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010011" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010100" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010101" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "1001100";
            
            when "0111010110" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111010111" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011000" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011001" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011010" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011011" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011100" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011101" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011110" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111011111" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "1001100";
            
            when "0111100000" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100001" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100010" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100011" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100100" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100101" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100110" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111100111" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111101000" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111101001" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "1001100";
            
            when "0111101010" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111101011" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111101100" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111101101" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111101110" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111101111" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111110000" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111110001" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111110010" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111110011" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "1001100";
            
            when "0111110100" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111110101" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111110110" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111110111" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111000" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111001" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111010" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111011" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111100" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111101" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0100100";
            
            when "0111111110" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "0111111111" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000000" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000001" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000010" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000011" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000100" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000101" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000110" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000000111" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0100100";
            
            when "1000001000" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001001" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001010" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001011" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001100" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001101" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001110" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000001111" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000010000" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000010001" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0100100";
            
            when "1000010010" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000010011" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000010100" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000010101" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000010110" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000010111" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000011000" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000011001" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000011010" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000011011" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0100100";
            
            when "1000011100" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000011101" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000011110" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000011111" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100000" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100001" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100010" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100011" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100100" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100101" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0100100";
            
            when "1000100110" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000100111" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101000" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101001" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101010" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101011" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101100" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101101" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101110" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000101111" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "0100100";
            
            when "1000110000" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110001" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110010" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110011" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110100" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110101" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110110" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000110111" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000111000" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000111001" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "0100100";
            
            when "1000111010" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1000111011" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1000111100" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1000111101" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1000111110" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1000111111" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1001000000" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1001000001" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1001000010" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1001000011" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "0100100";
            
            when "1001000100" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001000101" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001000110" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001000111" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001000" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001001" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001010" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001011" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001100" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001101" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "0100100";
            
            when "1001001110" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001001111" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010000" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010001" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010010" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010011" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010100" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010101" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010110" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when "1001010111" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0100100";
            
            when others =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0100100";
            end case;


            

    end process;
    
    
end behav ;